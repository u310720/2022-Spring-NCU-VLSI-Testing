`include "enum.sv"

module FSM (
    // Input
    input clk,
    input rst,
    
    // Output
    output logic [27:0] sel
);
    logic [4:0] cs, ns;

    always_ff @( posedge clk ) begin : CurrentState
        if (rst) begin
            cs <= FaultFree;
        end
        else begin
            cs <= ns;
        end
        // if (rst) begin
        //     cs <= FaultFree;
        // end
        // else begin
        //     if (cs == LoadAns) begin
        //         cs <= A_0;
        //     end
        //     else begin
        //         cs <= cs + 5'b1;
        //     end
        // end
    end

    always_comb begin : NextState
        if (cs == LoadAns) begin
            ns = A_0;
        end
        else begin
            ns = cs + 5'b1;
        end
    end

    always_comb begin : decoder
        case (cs)
            A_0: sel = 28'b0000_0000_0000_0000_0000_0000_0001;
            B_0: sel = 28'b0000_0000_0000_0000_0000_0000_0010;
            C_0: sel = 28'b0000_0000_0000_0000_0000_0000_0100;
            D_0: sel = 28'b0000_0000_0000_0000_0000_0000_1000;
            E_0: sel = 28'b0000_0000_0000_0000_0000_0001_0000;
            F_0: sel = 28'b0000_0000_0000_0000_0000_0010_0000;
            G_0: sel = 28'b0000_0000_0000_0000_0000_0100_0000;
            H_0: sel = 28'b0000_0000_0000_0000_0000_1000_0000;
            I_0: sel = 28'b0000_0000_0000_0000_0001_0000_0000;
            J_0: sel = 28'b0000_0000_0000_0000_0010_0000_0000;
            K_0: sel = 28'b0000_0000_0000_0000_0100_0000_0000;
            L_0: sel = 28'b0000_0000_0000_0000_1000_0000_0000;
            M_0: sel = 28'b0000_0000_0000_0001_0000_0000_0000;
            A_1: sel = 28'b0000_0000_0000_0010_0000_0000_0000;
            B_1: sel = 28'b0000_0000_0000_0100_0000_0000_0000;
            C_1: sel = 28'b0000_0000_0000_1000_0000_0000_0000;
            D_1: sel = 28'b0000_0000_0001_0000_0000_0000_0000;
            E_1: sel = 28'b0000_0000_0010_0000_0000_0000_0000;
            F_1: sel = 28'b0000_0000_0100_0000_0000_0000_0000;
            G_1: sel = 28'b0000_0000_1000_0000_0000_0000_0000;
            H_1: sel = 28'b0000_0001_0000_0000_0000_0000_0000;
            I_1: sel = 28'b0000_0010_0000_0000_0000_0000_0000;
            J_1: sel = 28'b0000_0100_0000_0000_0000_0000_0000;
            K_1: sel = 28'b0000_1000_0000_0000_0000_0000_0000;
            L_1: sel = 28'b0001_0000_0000_0000_0000_0000_0000;
            M_1: sel = 28'b0010_0000_0000_0000_0000_0000_0000;
            FaultFree: sel = 28'b0100_0000_0000_0000_0000_0000_0000;
            LoadAns: sel = 28'b1000_0000_0000_0000_0000_0000_0000;
            default: sel = 28'bxxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx;
        endcase
    end
endmodule