module SA0 (
    // Input
    input in,
    
    // Output
    output out
);
    assign out = 1'b0;
endmodule

module SA1 (
    // Input
    input in,
    
    // Output
    output out
);
    assign out = 1'b1;
endmodule