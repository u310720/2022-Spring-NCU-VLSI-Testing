`ifndef __ENUM_
`define __ENUM_
typedef enum logic [4:0] { 
    A_0, B_0, C_0, D_0, E_0, F_0, G_0, H_0, I_0, J_0, K_0, L_0, M_0,
    A_1, B_1, C_1, D_1, E_1, F_1, G_1, H_1, I_1, J_1, K_1, L_1, M_1, FaultFree, LoadAns
} faultlist;
`endif // __ENUM_